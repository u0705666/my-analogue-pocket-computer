module riscv_cpu(
    input clk,
    input reset_n
);

endmodule